module ULA(A, B, Reset, S);
	input [5:0] A, [5:0] B;
	input Reset;
	input [3:0] S;
	
	always @(*) begin
	// Implementar codigo
	end
endmodule